netcdf a {
dimensions:
        sample = 2304 ;
        z = 79 ;
variables:
        float latitude(sample) ;
                latitude:_FillValue = NaNf ;
                latitude:fortran_name = "\"xlat\"" ;
                latitude:standard_name = "\"latitude\"" ;
                latitude:long_name = "\"grid latitude in radians\"" ;
                latitude:field_dims = "\"(horizontal_dimension)\"" ;
                latitude:type = "\"real\"" ;
                latitude:kind = "\"kind_phys\"" ;
                latitude:intent = "\"in\"" ;
                latitude:optional = "\"F\"" ;
                latitude:units = "\"radians\"" ;
                latitude:coordinates = "tile time" ;
        float longitude(sample) ;
                longitude:_FillValue = NaNf ;
                longitude:fortran_name = "\"xlon\"" ;
                longitude:standard_name = "\"longitude\"" ;
                longitude:long_name = "\"grid longitude in radians\"" ;
                longitude:field_dims = "\"(horizontal_dimension)\"" ;
                longitude:type = "\"real\"" ;
                longitude:kind = "\"kind_phys\"" ;
                longitude:intent = "\"in\"" ;
                longitude:optional = "\"F\"" ;
                longitude:units = "\"radians\"" ;
                longitude:coordinates = "tile time" ;
        float pressure_thickness_of_atmospheric_layer(sample, z) ;
                pressure_thickness_of_atmospheric_layer:_FillValue = NaNf ;
                pressure_thickness_of_atmospheric_layer:standard_name = "\"air_pressure_difference_between_midlayers\"" ;
                pressure_thickness_of_atmospheric_layer:fortran_name = "\"del\"" ;
                pressure_thickness_of_atmospheric_layer:long_name = "\"pressure level thickness\"" ;
                pressure_thickness_of_atmospheric_layer:field_dims = "[\"horizontal_dimension\", \"vertical_dimension\"]" ;
                pressure_thickness_of_atmospheric_layer:type = "\"real\"" ;
                pressure_thickness_of_atmospheric_layer:kind = "\"kind_phys\"" ;
                pressure_thickness_of_atmospheric_layer:intent = "\"in\"" ;
                pressure_thickness_of_atmospheric_layer:optional = "\"F\"" ;
                pressure_thickness_of_atmospheric_layer:units = "\"Pa\"" ;
                pressure_thickness_of_atmospheric_layer:coordinates = "tile time" ;
        float air_pressure(sample, z) ;
                air_pressure:_FillValue = NaNf ;
                air_pressure:fortran_name = "\"prsl\"" ;
                air_pressure:standard_name = "\"air_pressure\"" ;
                air_pressure:long_name = "\"layer mean air pressure\"" ;
                air_pressure:field_dims = "[\"horizontal_dimension\", \"vertical_dimension\"]" ;
                air_pressure:type = "\"real\"" ;
                air_pressure:kind = "\"kind_phys\"" ;
                air_pressure:intent = "\"in\"" ;
                air_pressure:optional = "\"F\"" ;
                air_pressure:units = "\"Pa\"" ;
                air_pressure:coordinates = "tile time" ;
        float surface_air_pressure(sample) ;
                surface_air_pressure:_FillValue = NaNf ;
                surface_air_pressure:fortran_name = "\"ps\"" ;
                surface_air_pressure:standard_name = "\"surface_air_pressure\"" ;
                surface_air_pressure:long_name = "\"surface pressure\"" ;
                surface_air_pressure:field_dims = "[\"horizontal_dimension\"]" ;
                surface_air_pressure:type = "\"real\"" ;
                surface_air_pressure:kind = "\"kind_phys\"" ;
                surface_air_pressure:intent = "\"in\"" ;
                surface_air_pressure:optional = "\"F\"" ;
                surface_air_pressure:units = "\"Pa\"" ;
                surface_air_pressure:coordinates = "tile time" ;
        float air_temperature_input(sample, z) ;
                air_temperature_input:_FillValue = NaNf ;
                air_temperature_input:fortran_name = "\"t\"" ;
                air_temperature_input:standard_name = "\"air_temperature\"" ;
                air_temperature_input:long_name = "\"layer mean air temperature\"" ;
                air_temperature_input:field_dims = "[\"horizontal_dimension\", \"vertical_dimension\"]" ;
                air_temperature_input:type = "\"real\"" ;
                air_temperature_input:kind = "\"kind_phys\"" ;
                air_temperature_input:intent = "\"inout\"" ;
                air_temperature_input:optional = "\"F\"" ;
                air_temperature_input:units = "\"K\"" ;
                air_temperature_input:coordinates = "tile time" ;
        float specific_humidity_input(sample, z) ;
                specific_humidity_input:_FillValue = NaNf ;
                specific_humidity_input:fortran_name = "\"q\"" ;
                specific_humidity_input:standard_name = "\"specific_humidity\"" ;
                specific_humidity_input:long_name = "\"water vapor specific humidity\"" ;
                specific_humidity_input:field_dims = "[\"horizontal_dimension\", \"vertical_dimension\"]" ;
                specific_humidity_input:type = "\"real\"" ;
                specific_humidity_input:kind = "\"kind_phys\"" ;
                specific_humidity_input:intent = "\"inout\"" ;
                specific_humidity_input:optional = "\"F\"" ;
                specific_humidity_input:units = "\"kg kg-1\"" ;
                specific_humidity_input:coordinates = "tile time" ;
        float cloud_water_mixing_ratio_input(sample, z) ;
                cloud_water_mixing_ratio_input:_FillValue = NaNf ;
                cloud_water_mixing_ratio_input:fortran_name = "\"cwm\"" ;
                cloud_water_mixing_ratio_input:standard_name = "\"cloud_water_mixing_ratio\"" ;
                cloud_water_mixing_ratio_input:long_name = "\"moist cloud condensed water mixing ratio\"" ;
                cloud_water_mixing_ratio_input:field_dims = "[\"horizontal_dimension\", \"vertical_dimension\"]" ;
                cloud_water_mixing_ratio_input:type = "\"real\"" ;
                cloud_water_mixing_ratio_input:kind = "\"kind_phys\"" ;
                cloud_water_mixing_ratio_input:intent = "\"out\"" ;
                cloud_water_mixing_ratio_input:optional = "\"F\"" ;
                cloud_water_mixing_ratio_input:units = "\"kg kg-1\"" ;
                cloud_water_mixing_ratio_input:coordinates = "tile time" ;
        float air_temperature_after_last_gscond(sample, z) ;
                air_temperature_after_last_gscond:_FillValue = NaNf ;
                air_temperature_after_last_gscond:fortran_name = "\"tp\"" ;
                air_temperature_after_last_gscond:standard_name = "\"air_temperature_after_last_gscond\"" ;
                air_temperature_after_last_gscond:long_name = "\"air temperature after gscond was last called\"" ;
                air_temperature_after_last_gscond:field_dims = "[\"horizontal_dimension\", \"vertical_dimension\"]" ;
                air_temperature_after_last_gscond:type = "\"real\"" ;
                air_temperature_after_last_gscond:kind = "\"kind_phys\"" ;
                air_temperature_after_last_gscond:intent = "\"inout\"" ;
                air_temperature_after_last_gscond:optional = "\"F\"" ;
                air_temperature_after_last_gscond:units = "\"K\"" ;
                air_temperature_after_last_gscond:coordinates = "tile time" ;
        float specific_humidity_after_last_gscond(sample, z) ;
                specific_humidity_after_last_gscond:_FillValue = NaNf ;
                specific_humidity_after_last_gscond:fortran_name = "\"qp1\"" ;
                specific_humidity_after_last_gscond:standard_name = "\"specific_humidity_after_last_gscond\"" ;
                specific_humidity_after_last_gscond:long_name = "\"water vapor specific humidity after gscond was last called\"" ;
                specific_humidity_after_last_gscond:field_dims = "[\"horizontal_dimension\", \"vertical_dimension\"]" ;
                specific_humidity_after_last_gscond:type = "\"real\"" ;
                specific_humidity_after_last_gscond:kind = "\"kind_phys\"" ;
                specific_humidity_after_last_gscond:intent = "\"inout\"" ;
                specific_humidity_after_last_gscond:optional = "\"F\"" ;
                specific_humidity_after_last_gscond:units = "\"kg kg-1\"" ;
                specific_humidity_after_last_gscond:coordinates = "tile time" ;
        float surface_air_pressure_after_last_gscond(sample) ;
                surface_air_pressure_after_last_gscond:_FillValue = NaNf ;
                surface_air_pressure_after_last_gscond:fortran_name = "\"psp1\"" ;
                surface_air_pressure_after_last_gscond:standard_name = "\"surface_air_pressure_after_last_gscond\"" ;
                surface_air_pressure_after_last_gscond:long_name = "\"surface air surface pressure after gscond was last called\"" ;
                surface_air_pressure_after_last_gscond:field_dims = "[\"horizontal_dimension\"]" ;
                surface_air_pressure_after_last_gscond:type = "\"real\"" ;
                surface_air_pressure_after_last_gscond:kind = "\"kind_phys\"" ;
                surface_air_pressure_after_last_gscond:intent = "\"inout\"" ;
                surface_air_pressure_after_last_gscond:optional = "\"F\"" ;
                surface_air_pressure_after_last_gscond:units = "\"Pa\"" ;
                surface_air_pressure_after_last_gscond:coordinates = "tile time" ;
        float specific_humidity_after_gscond(sample, z) ;
                specific_humidity_after_gscond:_FillValue = NaNf ;
                specific_humidity_after_gscond:units = "unknown" ;
                specific_humidity_after_gscond:coordinates = "tile time" ;
        float air_temperature_after_gscond(sample, z) ;
                air_temperature_after_gscond:_FillValue = NaNf ;
                air_temperature_after_gscond:units = "unknown" ;
                air_temperature_after_gscond:coordinates = "tile time" ;
        float cloud_water_mixing_ratio_after_gscond(sample, z) ;
                cloud_water_mixing_ratio_after_gscond:_FillValue = NaNf ;
                cloud_water_mixing_ratio_after_gscond:units = "unknown" ;
                cloud_water_mixing_ratio_after_gscond:coordinates = "tile time" ;
        float air_temperature_after_precpd(sample, z) ;
                air_temperature_after_precpd:_FillValue = NaNf ;
                air_temperature_after_precpd:units = "unknown" ;
                air_temperature_after_precpd:coordinates = "tile time" ;
        float specific_humidity_after_precpd(sample, z) ;
                specific_humidity_after_precpd:_FillValue = NaNf ;
                specific_humidity_after_precpd:units = "unknown" ;
                specific_humidity_after_precpd:coordinates = "tile time" ;
        float cloud_water_mixing_ratio_after_precpd(sample, z) ;
                cloud_water_mixing_ratio_after_precpd:_FillValue = NaNf ;
                cloud_water_mixing_ratio_after_precpd:units = "unknown" ;
                cloud_water_mixing_ratio_after_precpd:coordinates = "tile time" ;
        float total_precipitation(sample) ;
                total_precipitation:_FillValue = NaNf ;
                total_precipitation:fortran_name = "\"rn\"" ;
                total_precipitation:standard_name = "\"total_precipitation\"" ;
                total_precipitation:long_name = "\"explicit precipitation amount on physics timestep\"" ;
                total_precipitation:field_dims = "[\"horizontal_dimension\"]" ;
                total_precipitation:type = "\"real\"" ;
                total_precipitation:kind = "\"kind_phys\"" ;
                total_precipitation:intent = "\"out\"" ;
                total_precipitation:optional = "\"F\"" ;
                total_precipitation:units = "\"m\"" ;
                total_precipitation:coordinates = "tile time" ;
        float ratio_of_snowfall_to_rainfall(sample) ;
                ratio_of_snowfall_to_rainfall:_FillValue = NaNf ;
                ratio_of_snowfall_to_rainfall:fortran_name = "\"sr\"" ;
                ratio_of_snowfall_to_rainfall:standard_name = "\"ratio_of_snowfall_to_rainfall\"" ;
                ratio_of_snowfall_to_rainfall:long_name = "\"ratio of snowfall to large-scale rainfall\"" ;
                ratio_of_snowfall_to_rainfall:field_dims = "[\"horizontal_dimension\"]" ;
                ratio_of_snowfall_to_rainfall:type = "\"real\"" ;
                ratio_of_snowfall_to_rainfall:kind = "\"kind_phys\"" ;
                ratio_of_snowfall_to_rainfall:intent = "\"out\"" ;
                ratio_of_snowfall_to_rainfall:optional = "\"F\"" ;
                ratio_of_snowfall_to_rainfall:units = "\"frac\"" ;
                ratio_of_snowfall_to_rainfall:coordinates = "tile time" ;
        float tendency_of_rain_water_mixing_ratio_due_to_microphysics(sample, z) ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:_FillValue = NaNf ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:fortran_name = "\"rainp\"" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:standard_name = "\"tendency_of_rain_water_mixing_ratio_due_to_microphysics\"" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:long_name = "\"tendency of rain water mixing ratio due to microphysics\"" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:field_dims = "[\"horizontal_dimension\", \"vertical_dimension\"]" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:type = "\"real\"" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:kind = "\"kind_phys\"" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:intent = "\"out\"" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:optional = "\"F\"" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:units = "\"kg kg-1 s-1\"" ;
                tendency_of_rain_water_mixing_ratio_due_to_microphysics:coordinates = "tile time" ;
        int64 time ;
                time:units = "days since 2016-04-25 03:45:00.000000" ;
                time:calendar = "julian" ;
        int64 tile ;
}